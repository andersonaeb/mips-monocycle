----------------------------------------------------------------------------------
-- MIPS MONOCYCLE
-- Datapath 
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MixMonocycle is
	
end MixMonocycle;

-------------------------------------------------------------------------

architecture behavior of MixMonocycle is
	

	
begin
	
end behavior;